LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY LED7S IS
PORT(  CLK : IN STD_LOGIC;
         D0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 D1: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 D2: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 D3: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 
		 EN: IN STD_LOGIC;
		  C: BUFFER STD_LOGIC_VECTOR(2 DOWNTO 0);
	 LED7S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END;

ARCHITECTURE ONE OF LED7S IS
  SIGNAL D: STD_LOGIC_VECTOR(3 DOWNTO 0);
 
BEGIN


P1:PROCESS(CLK, EN)
BEGIN 
	IF CLK'EVENT AND CLK='1' THEN
		IF C < "011" THEN 
			C <= C+1;
		ELSE
			C<="000";
		END IF;
	END IF;
	
IF EN = '0' THEN
	IF CLK'EVENT AND CLK='1' THEN
		IF D < "1111" THEN
			D <= D + 1;
		ELSE
			D <= "0000";
		END IF;
	END IF;
ELSE
	IF C = "000" THEN
		D <= D0;
	END IF;
	IF C = "001" THEN
		D <= D1;
	END IF;
	IF C = "010" THEN
		D <= D2;
	END IF;
	IF C = "011" THEN
		D <= D3;
	END IF;
END IF;
END PROCESS P1;

P2:PROCESS(D)
BEGIN
 CASE D IS
 WHEN"0000"=>LED7S<="00111111";
 WHEN"0001"=>LED7S<="00000110";
 WHEN"0010"=>LED7S<="01011011";
 WHEN"0011"=>LED7S<="01001111";
 WHEN"0100"=>LED7S<="01100110";
 WHEN"0101"=>LED7S<="01101101";
 WHEN"0110"=>LED7S<="01111101";
 WHEN"0111"=>LED7S<="00000111";
 WHEN"1000"=>LED7S<="01111111";
 WHEN"1001"=>LED7S<="01101111";
 WHEN"1010"=>LED7S<="01110111";
 WHEN"1011"=>LED7S<="01111100";
 WHEN"1100"=>LED7S<="00111001";
 WHEN"1101"=>LED7S<="01011110";
 WHEN"1110"=>LED7S<="01111001";
 WHEN"1111"=>LED7S<="01110001";
 WHEN OTHERS=>NULL;
 END CASE;
 END PROCESS P2; 
 
 
       
END ONE;
	